// Test Verilog module
module mac (
    output     reg[0:15] out,
    input       reg[0:15] ina, inb, 
    input       clk, sclrn
);



endmodule
